`include "defines.v"

module exu_oitf(
    output                  dis_ready,

    input                   dis_ena,
    input                   ret_ena

    // output  [`ITAG]
);

endmodule
